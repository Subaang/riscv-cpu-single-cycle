module top (
    input clk,
    input reset
);

    // Instantiate modules (PC, RegFile, ALU, etc.) here later

endmodule
