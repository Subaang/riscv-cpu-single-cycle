module Top (
    input logic clk,
    input logic reset
);

    // Instantiate modules (PC, RegFile, ALU, etc.) here later

endmodule
